library IEEE;
use IEEE.std_logic_1164.ALL;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use work.vga_controller_cfg.all;

--safe implementation yes
architecture tools_arch of tlv_pc_ifc is

  signal vga_mode: std_logic_vector(60 downto 0);
  signal red: std_logic_vector(2 downto 0);
  signal green: std_logic_vector(2 downto 0);
  signal blue: std_logic_vector(2 downto 0);
  signal rgb : std_logic_vector(8 downto 0);

  signal vgaRow: std_logic_vector(11 downto 0);
  signal vgaCol: std_logic_vector(11 downto 0);

  signal keyboard	: std_logic_vector(15 downto 0);

  signal fps: std_logic;
	
  type six is 
  record
	r : std_logic_vector(1 downto 0);
	g : std_logic_vector(1 downto 0);
	b : std_logic_vector(1 downto 0);
  end record;
  
  type nine is
  record
	r : std_logic_vector(2 downto 0);
	g : std_logic_vector(2 downto 0);
	b : std_logic_vector(2 downto 0);
  end record;
  
  signal bgColor: six := ("00", "00", "00");
  
  --lets have 16 colors
  type pallete is array (0 to 15) of nine;
  constant colorPallete : pallete := (
	0 => ("000", "000", "000"),
	1 => ("101", "000", "000"),
	2 => ("110", "000", "000"),
	3 => ("111", "000", "000"),
	others => ("000", "000", "000")
  );
  
  function repairPos(input : integer) return integer is
  variable result : integer range 0 to 14;
  begin
	if(input > 14) then
		result := 14;
	else
		result := input;
	end if;
	return result;
  end function;
  
  function pallete2color(input : std_logic_vector(1 downto 0)) return nine is
  variable result : nine;
  begin
    case input is
		when "00" =>
			result := colorPallete(0); 
		when "01" =>
			result := colorPallete(1);
		when "10" =>
			result := colorPallete(2);
		when "11" =>
			result := colorPallete(3);
		when others =>
			result := colorPallete(0);
	 end case;
	 return result;
  end function;
  
  function color2nine(input : nine) return std_logic_vector is
  variable tmp : std_logic_vector(8 downto 0);
  begin
   tmp := input.r & input.g & input.b;
	return tmp;
  end function;
  
  function letterBitmap(input : character) return integer is
  variable result : integer range 1 to 27;
  begin
    case input is
		when 'A' =>
			result := 1;
		when 'B' =>
			result := 2;
		when 'C' =>
			result := 3;
		when 'D' =>
			result := 4;
		when 'E' =>
			result := 5;
		when 'F' =>
			result := 6;
		when 'G' =>
			result := 7;
		when 'H' =>
			result := 8;
		when 'I' =>
			result := 9;
		when 'J' =>
			result := 10;
		when 'K' =>
			result := 11;
		when 'L' =>
			result := 12;
		when 'M' =>
			result := 13;
		when 'N' =>
			result := 14;
		when 'O' =>
			result := 15;
		when 'P' =>
			result := 16;
		when 'Q' =>
			result := 17;
		when 'R' =>
			result := 18;
		when 'S' =>
			result := 19;
		when 'T' =>
			result := 20;
		when 'U' =>
			result := 21;
		when 'V' =>
			result := 22;
		when 'W' =>
			result := 23;
		when 'X' =>
			result := 24;
		when 'Y' =>
			result := 25;
		when 'Z' =>
			result := 26;
		when ' ' =>
			result := 27;
		when others => result := 27;
	end case;
	return result;
  end function;
  
  --to store bitmap of single letters
  --type bitmap_row is array (0 to 14) of std_logic_vector(1 downto 0);
  --type bitmap is array(0 to 14) of bitmap_row;
  
  type bitmap2 is array(0 to 224) of std_logic_vector(1 downto 0);
  
  constant LETTER_SIZE : integer := 14;
  
  type letter_entity is
  record
    x : std_logic_vector(9 downto 0);
	 y : std_logic_vector(9 downto 0);
    c : character;
  end record;	 
  constant END_LETTER : letter_entity := (
    x => "0000000000",
	 y => "0000000000",
	 c => ' '
  );
  
  --number of letter entities (letters to draw)
  constant num_entities : integer := 5;
  
  type list is array (1 to num_entities) of letter_entity;
  
  signal entity_list : list := ( others => (x => "0000000000", y => "0000000000", c => ' '));
  
  type letter_list is array (1 to 26) of bitmap2;
  
  signal letter_rom : letter_list := (
  1 => (
    --A
			"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"11", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", "01", "10", "10", "10"
  ),	
	2 => (
    --B
			"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"11", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", "00", 
			"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "01", "00", "00", "10", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
	),
	3 => (
    --C
			"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", 
			"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "01", "10", "10", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
			"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
	),
4 => (
    --D
			"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
	),		
5 => (
    --E
			"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", 
			"11", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "01", "10", "10", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "01", "11", "11", "11", "11", "11", "01", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", 
			"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
			"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
	),		
6 => (
    --F
			"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", 
			"11", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "01", "10", "10", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", 
			"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00"
	 ),
7 => (
    --G
			"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", 
			"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "01", "10", "10", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "11", "11", "11", "11", "11", "01", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "01", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
	 ),
8 => (
    --H
			"11", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
			"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
			"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
			"01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", "01", "10", "10", "10"
	 ),
9 => (
		--I
				"00", "00", "00", "00", "11", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", 
				"00", "00", "00", "00", "01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00" 
), 
10 => (
		--J
				"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "01", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
				"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "11", "11", "11", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
),
11 => (
		--K
				"11", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", "00", 
				"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", "01", "10", "10", "10"
), 
12 => (
		--L
				"11", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
				"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
), 
13 => (
		--M
				"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"11", "00", "00", "01", "10", "10", "10", "01", "00", "10", "10", "01", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "01", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "11", "00", "10", "00", "11", "00", "00", "10", 
				"01", "10", "10", "10", "10", "10", "00", "01", "10", "10", "00", "01", "10", "10", "10"
), 
14 => (
		--N
				"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", "01", "10", "10", "10"
), 
15 => (
		--O
				"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
), 
16 => (
		--P
				"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"11", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00"
), 
17 => (
		--Q
				"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "00", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", "00", "00", 
				"11", "00", "00", "01", "10", "10", "10", "10", "10", "01", "00", "00", "10", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", "00", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", "00", "00", 
				"11", "00", "00", "01", "11", "01", "00", "00", "00", "11", "00", "00", "10", "00", "00", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "01", "10", "10", "10", "00", "00", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "01", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10"
), 
18 => (
--R
"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", "00", 
"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", "01", "10", "10", "10"
), 
19 => (
--S
"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", 
"11", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "01", "10", "10", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "11", "11", "11", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"

), 
20 => (
--T
"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", 
"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "01", 
"11", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "01", "10", "10", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
"01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00"
), 
21 => (
--U
"11", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
"00", "01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
), 
22 => (
--V
"11", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"01", "00", "00", "01", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"00", "10", "00", "00", "11", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
"00", "00", "10", "00", "00", "11", "11", "11", "00", "00", "00", "11", "00", "00", "10", 
"00", "00", "00", "10", "00", "00", "00", "00", "11", "00", "00", "11", "00", "00", "10", 
"00", "00", "00", "00", "10", "00", "00", "00", "00", "11", "00", "11", "00", "00", "10", 
"00", "00", "00", "00", "00", "10", "00", "00", "00", "00", "11", "11", "00", "00", "10", 
"00", "00", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "10", 
"00", "00", "00", "00", "00", "00", "00", "10", "10", "10", "10", "10", "10", "10", "00"
), 
23 => (
		--W
				"11", "11", "11", "01", "00", "00", "11", "11", "01", "00", "00", "11", "11", "11", "01", 
				"11", "00", "00", "10", "00", "00", "11", "00", "10", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "11", "00", "10", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "11", "00", "10", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "11", "00", "10", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "11", "00", "10", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "01", "10", "10", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"00", "01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
), 
24 => (
		--X
				"11", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"00", "11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", "00", 
				"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"01", "10", "10", "10", "10", "10", "00", "00", "00", "00", "00", "01", "10", "10", "10"
), 
25 => (
		--Y
				"11", "11", "11", "01", "00", "00", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "01", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
				"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "11", "11", "11", "11", "01", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"00", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00"
		
), 
26 => (
		--Z
				"11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "01", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"11", "00", "00", "10", "10", "10", "10", "10", "10", "10", "10", "01", "00", "00", "10", 
				"01", "10", "10", "10", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"00", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"11", "00", "00", "01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "00", 
				"11", "00", "00", "10", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", 
				"11", "00", "00", "01", "11", "01", "00", "00", "00", "00", "00", "11", "11", "11", "01", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "10", "00", "00", "00", "00", "00", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "01", "11", "11", "11", "11", "11", "11", "00", "00", "10", 
				"11", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "00", "10", 
				"01", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10", "10"
)
  );
  
  --drawing functions / procedures
--convert function from 2-2-2 rgb to 3-3-3
function RGB_6to9(input : six) return std_logic_vector is
	variable tmp : std_logic_vector(8 downto 0); 
begin
	if(input.r = 0) then
		tmp(8 downto 6) := "000";
	else
		tmp(8 downto 7) := input.r;
		tmp(6) := '1';
	end if;
	
	if(input.g = 0) then
		tmp(5 downto 3) := "000";
	else
		tmp(5 downto 4) := input.g;
		tmp(3) := '1';
	end if;
	
	if(input.b = 0) then
		tmp(2 downto 0) := "000";
	else
		tmp(2 downto 1) := input.b;
		tmp(0) := '1';
	end if;
	
	return tmp;
end function;

component keyboard_controller
	port(
		CLK      : in std_logic;
		RST      : in std_logic;
		
		DATA_OUT : out std_logic_vector(15 downto 0);
		DATA_VLD : out std_logic;
		
		KB_KIN   : out std_logic_vector(3 downto 0);
		KB_KOUT  : in  std_logic_vector(3 downto 0)
	);
end component;

begin

kbrd_ctrl: entity work.keyboard_controller(arch_keyboard)
port map (
	CLK => CLK,
	RST => RESET,
	
	DATA_OUT => keyboard,
	DATA_VLD => open,
	
	KB_KIN   => KIN,
	KB_KOUT  => KOUT
);


fps_generator: entity work.engen generic map ( MAXVALUE => 9000000) port map ( CLK => CLK, ENABLE => '1', EN => fps );

vga: entity work.vga_controller(arch_vga_controller)
  port map(
    CLK => CLK,
    RST => RESET,
    ENABLE => '1',
    MODE => vga_mode,
    DATA_RED => red,
    DATA_GREEN => green,
    DATA_BLUE => blue,
    ADDR_COLUMN => vgaCol,
    ADDR_ROW => vgaRow,
    VGA_RED => RED_V,
    VGA_GREEN => GREEN_V,
    VGA_BLUE => BLUE_V,
    VGA_HSYNC => HSYNC_V,
    VGA_VSYNC => VSYNC_V
  );
  
setmode(r640x480x60, vga_mode);

-- user code here!
app_logic: process(fps)
	variable cursor_x : integer;
	variable cursor_y : integer;
	variable latch : bit := '0';
	variable init : bit := '1';
	variable divider : bit := '0';
begin
	if(fps'event and fps = '1') then
		if(init = '1')then
			cursor_x := 280;
			cursor_y := 225;
			entity_list(1).x <= std_logic_vector(to_unsigned(cursor_x, 10));
			entity_list(1).y <= std_logic_vector(to_unsigned(cursor_y, 10));
			entity_list(1).c <= 'H';
			cursor_x := cursor_x + LETTER_SIZE;
			entity_list(2).x <= std_logic_vector(to_unsigned(cursor_x, 10));
			entity_list(2).y <= std_logic_vector(to_unsigned(cursor_y, 10));
			entity_list(2).c <= 'E';
			cursor_x := cursor_x + LETTER_SIZE;
			entity_list(3).x <= std_logic_vector(to_unsigned(cursor_x, 10));
			entity_list(3).y <= std_logic_vector(to_unsigned(cursor_y, 10));
			entity_list(3).c <= 'L';
			cursor_x := cursor_x + LETTER_SIZE;
			entity_list(4).x <= std_logic_vector(to_unsigned(cursor_x, 10));
			entity_list(4).y <= std_logic_vector(to_unsigned(cursor_y, 10));
			entity_list(4).c <= 'L';
			cursor_x := cursor_x + LETTER_SIZE;
			entity_list(5).x <= std_logic_vector(to_unsigned(cursor_x, 10));
			entity_list(5).y <= std_logic_vector(to_unsigned(cursor_y, 10));
			entity_list(5).c <= 'O';
			init := '0';
		end if;
		if(divider = '1') then
			if(latch = '0') then
				entity_list(1).c <= 'H';
				entity_list(2).c <= 'E';
				entity_list(3).c <= 'L';
				entity_list(4).c <= 'L';
				entity_list(5).c <= 'O';
				latch := '1';
			else
				entity_list(1).c <= 'W';
				entity_list(2).c <= 'O';
				entity_list(3).c <= 'R';
				entity_list(4).c <= 'L';
				entity_list(5).c <= 'D';
				latch := '0';
			end if;
			divider := '0';
		else
			divider := '1';
		end if;
	end if;
end process;

-- DO NOT CHANGE THIS
draw: process(CLK)
	variable pos_x : integer range 0 to 14;
	variable pos_y  : integer range 0 to 14;
	variable pos_c : integer range 0 to 224;
	variable letter_number : integer range 1 to 27;
	variable tmp_vector : std_logic_vector(1 downto 0);
	variable tmp_nine : nine;
	variable tmp_letter : bitmap2;
begin
	if(CLK'event and CLK = '1') then
		if(vgaRow < 479 and vgaCol < 639) then
				rgb <= RGB_6to9(bgColor);
				for i_object in 1 to num_entities loop
					if(entity_list(i_object) = END_LETTER) then
						exit;
					end if;
					
					if(vgaCol >= entity_list(i_object).x and vgaCol <= (entity_list(i_object).x + LETTER_SIZE)) then					
						if(vgaRow >= entity_list(i_object).y and vgaRow <= (entity_list(i_object).y + LETTER_SIZE)) then	
							pos_x := repairPos(conv_integer(vgaCol(9 downto 0) - entity_list(i_object).x));
							pos_y := repairPos(conv_integer(vgaRow(9 downto 0) - entity_list(i_object).y));
							letter_number := letterBitmap(entity_list(i_object).c);
							tmp_letter := letter_rom(letter_number);
							pos_c := pos_x + (pos_y * 15);
							tmp_vector := tmp_letter(pos_c);
							rgb <= color2nine(pallete2color(tmp_vector));
						end if;
					end if;
				end loop;
		else
			rgb <= RGB_6to9(bgColor);
		end if;

	end if;
end process;

red <= rgb(8 downto 6);
green <= rgb(5 downto 3);
blue <= rgb(2 downto 0);

end tools_arch;
